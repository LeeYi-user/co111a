module Nand(input a, b, output out);
    nand g(out, a, b);
endmodule
